library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use work.mario_package.all;

package vga_package is

	--types definition
	
	--MATRICE USATA DALLA FUNZIONE GET_COLOR PER RESTITUIRE LE 3 COMPONENTI RGB A 4 BIT
	type matrix_color is array (0 to 2) of std_logic_vector(3 downto 0);
	
	--CONSTANTS
	
	--game
	constant JUMP_UNIT						: positive := 125;
	
	constant GAME_WIDTH						: natural := 640;
	constant GAME_HEIGHT						: natural := 480;
		
	--VITE
	constant MAX_LIVES						: positive := 3;
	
	--bounds
	constant BOUND_TOP_THICKNESS			: natural := 50;
	constant BOUND_LAT_THICKNESS			: natural := 20;
	constant BOUND_TOP						: natural := BOUND_TOP_THICKNESS;
	constant BOUND_LEFT						: natural := BOUND_LAT_THICKNESS;
	constant BOUND_RIGHT						: natural := GAME_WIDTH-BOUND_LAT_THICKNESS;
	constant BOUND_BOTTOM					: natural := GAME_HEIGHT-16;
	
	--STARS LIFE
	constant STAR1_X 						: natural := 35;
	constant STAR1_Y 						: natural := 10;
	
	constant STAR2_X 						: natural := 70;
	constant STAR2_Y 						: natural := 10;
	
	constant STAR3_X 						: natural := 105;
	constant STAR3_Y 						: natural := 10;
	
	--TIMER IN PLAYING
	constant PRIMA_CIFRA_X 				: natural := 300;
	constant PRIMA_CIFRA_Y 				: natural := 10;
	
	constant SECONDA_CIFRA_X 			: natural := 320;
	constant SECONDA_CIFRA_Y 			: natural := 10;
	
	--PAUSE
	constant PAUSE_X 						: natural := 300;
	constant PAUSE_Y 						: natural := 10;
	
	--COIN SCORE
	constant COIN_SCORE_X 				: natural := 496;
	constant COIN_SCORE_Y 				: natural := 10;
	
	--X SCORE
	constant X_SCORE_X 				: natural := 514;
	constant X_SCORE_Y 				: natural := 10;
	
	--NUM COINS TO CATCH
	constant COIN_TO_CATCH_FIRST_X 				: natural := 532;
	constant COIN_TO_CATCH_FIRST_Y 				: natural := 10;
	
	constant COIN_TO_CATCH_SECOND_X 				: natural := 550;
	constant COIN_TO_CATCH_SECOND_Y 				: natural := 10;
	
	-- =
	constant EQUAL_X 				: natural := 568;
	constant EQUAL_Y 				: natural := 10;
	
	--MY SCORE
	constant MY_FIRST_SCORE_X 				: natural := 586;
	constant MY_FIRST_SCORE_Y 				: natural := 10;
	
	constant MY_SECOND_SCORE_X 				: natural := 604;
	constant MY_SECOND_SCORE_Y 				: natural := 10;
	
	--CLOUDS POSITION
	constant NUM_CLOUDS : natural := 6;
	
	constant CLOUD_1 : coord :=(
		x => 90,
		y => 200
	);
	constant CLOUD_2 : coord :=(
		x => 150,
		y => 90
	);
	constant CLOUD_3 : coord :=(
		x => 250,
		y => 150
	);
	constant CLOUD_4 : coord :=(
		x => 330,
		y => 300
	);	
	constant CLOUD_5 : coord :=(
		x => 448,
		y => 200
	);	
	constant CLOUD_6 : coord :=(
		x => 520,
		y => 330
	);	
	
	type t_clouds_array is array(0 to NUM_CLOUDS-1) of coord; -- coordinate type
	constant CLOUDS : t_clouds_array := (CLOUD_1, CLOUD_2, CLOUD_3, CLOUD_4, CLOUD_5, CLOUD_6); -- all the blocks are stored here
	
	--HILL POSITION
	constant HILL1_X 							: natural := 200;
	constant HILL1_Y 							: natural := 424;
	
	constant HILL2_X 							: natural := 500;
	constant HILL2_Y 							: natural := 424;
	
	--FLOOR POSITION
	constant FLOOR_X 							: natural := 20;
	constant FLOOR_Y 							: natural := 462;
	
	--BRICK POSITION
	constant BRICK_X 							: natural := 150;
	constant BRICK_Y 							: natural := 370;
	
	constant MARIO_STARTING_POSX			: natural := GAME_WIDTH/2-MARIO_WIDTH;
	constant MARIO_STARTING_POSY			: natural := 340;
	
	--screen
	constant VISIBLE_WIDTH    : natural := 640;
	constant VISIBLE_HEIGHT   : natural := 480;

	--vertical sync
	constant VERTICAL_FRONT_PORCH : natural := 10;
	constant VERTICAL_SYNC_PULSE : natural := 2;
	constant VERTICAL_BACK_PORCH : natural := 33;

	--horizontal sync
	constant HORIZONTAL_FRONT_PORCH : natural := 16;
	constant HORIZONTAL_SYNC_PULSE : natural := 96;
	constant HORIZONTAL_BACK_PORCH : natural := 48;
	
	--VGA screen
	constant TOTAL_W: integer := HORIZONTAL_FRONT_PORCH + HORIZONTAL_SYNC_PULSE +HORIZONTAL_BACK_PORCH + VISIBLE_WIDTH;	--800
	constant TOTAL_H: integer := VERTICAL_FRONT_PORCH + VERTICAL_SYNC_PULSE +VERTICAL_BACK_PORCH + VISIBLE_HEIGHT; --525

	constant WINDOW_HORIZONTAL_START: integer := HORIZONTAL_FRONT_PORCH + HORIZONTAL_SYNC_PULSE + HORIZONTAL_BACK_PORCH; 
	constant WINDOW_VERTICAL_START: integer := VERTICAL_FRONT_PORCH + VERTICAL_SYNC_PULSE +VERTICAL_BACK_PORCH;
	
		
	--MATRICE CHE MI INDICA SE IL PIXEL IDENTIFICA UN ELEMENTO DI MARIO
	type mario_form is array (0 to MARIO_HEIGHT - 1 , 0 to MARIO_WIDTH - 1) of std_logic;
	constant mario_borders : mario_form := (
	
		("0000001111100000"),
		("0000111111100000"),
		("0001111111100000"),
		("0001111111111100"),
		("0001111111110000"),
		("0011111111111100"),
		("0011111111111110"),
		("0111111111111110"),
		("0111111111111100"),
		("0111111111111100"),
		("0001111111111000"),
		("0000111111100000"),
		("0000111111110000"),
		("0001111111111000"),
		("0011111111111100"),
		("0111111111111110"),
		("0111111111111110"),
		("1111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("0111111111111110"),
		("0111111111111110"),
		("0011111111111100"),
		("0111111001111110"),
		("0111110000111110"),
		("0111110000111110"),
		("0011110000111100"),
		("0011110000111100"),
		("1111110000111111"),
		("1111110000111111")
	);	
	
	--MATRICE CHE RESTITUISCE IL COLORE DI OGNI PIXEL ASSOCIATO A MARIO
	type mario_colori is array (0 to MARIO_HEIGHT - 1 , 0 to MARIO_WIDTH - 1) of std_logic_vector(3 downto 0);
	constant mario_colors : mario_colori := (
		( x"0", x"0", x"0",  x"0",  x"0",  x"0",  x"2", x"2",  x"2",  x"2",  x"2", x"0",  x"0",  x"0", x"0",  x"0"),
		( x"0", x"0", x"0",  x"0",  x"2",  x"2",  x"2", x"2",  x"2",  x"2",  x"4", x"0",  x"0",  x"0", x"0",  x"0"),
		( x"0", x"0", x"0",  x"2",  x"2",  x"2",  x"2", x"2",  x"4",  x"4",  x"4", x"0",  x"0",  x"0", x"0",  x"0"),
		( x"0", x"0", x"0",  x"2",  x"2",  x"2",  x"2", x"2",  x"2",  x"2",  x"2", x"2",  x"2",  x"2", x"0",  x"0"),
		( x"0", x"0", x"0",  x"3",  x"3",  x"3",  x"1", x"1",  x"3",  x"1",  x"1", x"1",  x"0",  x"0", x"0",  x"0"),
		( x"0", x"0", x"3",  x"1",  x"1",  x"3",  x"1", x"1",  x"3",  x"3",  x"1", x"1",  x"1",  x"1", x"0",  x"0"),
		( x"0", x"0", x"3",  x"1",  x"1",  x"3",  x"3", x"1",  x"1",  x"1",  x"1", x"1",  x"1",  x"1", x"1",  x"0"),
		( x"0", x"3", x"3",  x"1",  x"1",  x"3",  x"3", x"1",  x"1",  x"1",  x"3", x"1",  x"1",  x"1", x"1",  x"0"),
		( x"0", x"3", x"3",  x"1",  x"1",  x"1",  x"1", x"1",  x"3",  x"3",  x"3", x"3",  x"3",  x"3", x"0",  x"0"),
		( x"0", x"3", x"3",  x"3",  x"1",  x"1",  x"1", x"1",  x"1",  x"3",  x"3", x"3",  x"3",  x"3", x"0",  x"0"),
		( x"0", x"0", x"0",  x"3",  x"3",  x"1",  x"1", x"1",  x"1",  x"1",  x"1", x"1",  x"1",  x"0", x"0",  x"0"),
		( x"0", x"0", x"0",  x"0",  x"2",  x"1",  x"1", x"1",  x"1",  x"1",  x"3", x"0",  x"0",  x"0", x"0",  x"0"),
		( x"0", x"0", x"0",  x"0",  x"3",  x"2",  x"3", x"3",  x"3",  x"3",  x"2", x"3",  x"0",  x"0", x"0",  x"0"),
		( x"0", x"0", x"0",  x"3",  x"3",  x"2",  x"3", x"3",  x"3",  x"3",  x"2", x"3",  x"3",  x"0", x"0",  x"0"),
		( x"0", x"0", x"3",  x"3",  x"3",  x"2",  x"3", x"3",  x"3",  x"3",  x"2", x"3",  x"3",  x"3", x"0",  x"0"),
		( x"0", x"3", x"3",  x"3",  x"3",  x"2",  x"3", x"3",  x"3",  x"3",  x"2", x"3",  x"3",  x"3", x"3",  x"0"),
		( x"0", x"3", x"3",  x"3",  x"2",  x"2",  x"3", x"3",  x"3",  x"3",  x"2", x"2",  x"3",  x"3", x"3",  x"0"),
		( x"3", x"3", x"3",  x"3",  x"2",  x"2",  x"3", x"3",  x"3",  x"3",  x"2", x"2",  x"3",  x"3", x"3",  x"3"),
		( x"3", x"3", x"3",  x"3",  x"2",  x"2",  x"2", x"2",  x"2",  x"2",  x"2", x"2",  x"3",  x"3", x"3",  x"3"),
		( x"3", x"3", x"3",  x"3",  x"2",  x"4",  x"2", x"2",  x"2",  x"2",  x"4", x"2",  x"3",  x"3", x"3",  x"3"),
		( x"1", x"1", x"1",  x"1",  x"2",  x"2",  x"2", x"2",  x"2",  x"2",  x"2", x"2",  x"1",  x"1", x"1",  x"1"),
		( x"1", x"1", x"1",  x"1",  x"2",  x"2",  x"2", x"2",  x"2",  x"2",  x"2", x"2",  x"1",  x"1", x"1",  x"1"),
		( x"0", x"1", x"1",  x"1",  x"2",  x"2",  x"2", x"2",  x"2",  x"2",  x"2", x"2",  x"1",  x"1", x"1",  x"0"),
		( x"0", x"1", x"1",  x"2",  x"2",  x"2",  x"2", x"2",  x"2",  x"2",  x"2", x"2",  x"2",  x"1", x"1",  x"0"),
		( x"0", x"0", x"2",  x"2",  x"2",  x"2",  x"2", x"2",  x"2",  x"2",  x"2", x"2",  x"2",  x"2", x"0",  x"0"),
		( x"0", x"2", x"2",  x"2",  x"2",  x"2",  x"2", x"0",  x"0",  x"2",  x"2", x"2",  x"2",  x"2", x"2",  x"0"),
		( x"0", x"2", x"2",  x"2",  x"2",  x"2",  x"0", x"0",  x"0",  x"0",  x"2", x"2",  x"2",  x"2", x"2",  x"0"),
		( x"0", x"2", x"2",  x"2",  x"2",  x"2",  x"0", x"0",  x"0",  x"0",  x"2", x"2",  x"2",  x"2", x"2",  x"0"),
		( x"0", x"0", x"3",  x"3",  x"3",  x"3",  x"0", x"0",  x"0",  x"0",  x"3", x"3",  x"3",  x"3", x"0",  x"0"),
		( x"0", x"0", x"3",  x"3",  x"3",  x"3",  x"0", x"0",  x"0",  x"0",  x"3", x"3",  x"3",  x"3", x"0",  x"0"),
		( x"3", x"3", x"3",  x"3",  x"3",  x"3",  x"0", x"0",  x"0",  x"0",  x"3", x"3",  x"3",  x"3", x"3",  x"3"),
		( x"3", x"3", x"3",  x"3",  x"3",  x"3",  x"0", x"0",  x"0",  x"0",  x"3", x"3",  x"3",  x"3", x"3",  x"3")
	);
	
	
	type cloud_form is array (0 to CLOUD_HEIGHT - 1 , 0 to CLOUD_WIDTH - 1) of std_logic;
	constant cloud_borders : cloud_form := (
		("0000000000000000000000000000111111110000000000000000000000000000"),
		("0000000000000000000000000000111111110000000000000000000000000000"),
		("0000000000000000000000000011111111111100000000000000000000000000"),
		("0000000000000000000000000011111111111100000000000000000000000000"),
		("0000000000000000000000111111111111111111000000000000000000000000"),
		("0000000000000000000000111111111111111111000000000000000000000000"),
		("0000000000000000000011111111111111111111111110000000000000000000"),
		("0000000000000000000011111111111111111111111110000000000000000000"),
		("0000000000000000000011111111111111111111111111100000000000000000"),
		("0000000000000000000011111111111111111111111111100000000000000000"),
		("0000000000000000000011111111111111111111111111110000000000000000"),
		("0000000000000000000011111111111111111111111111110000000000000000"),
		("0000000000000000001111111111111111111111111111110000000000000000"),
		("0000000000000000001111111111111111111111111111110000000000000000"),
		("0000000000000000111111111111111111111111111111110000000000000000"),
		("0000000000000000111111111111111111111111111111111111111100000000"),
		("0000000000111111111111111111111111111111111111111111111100000000"),
		("0000000000111111111111111111111111111111111111111111111111000000"),
		("0000000011111111111111111111111111111111111111111111111111000000"),
		("0000000011111111111111111111111111111111111111111111111111000000"),
		("0000001111111111111111111111111111111111111111111111111111000000"),
		("0000001111111111111111111111111111111111111111111111111111111100"),
		("0000011111111111111111111111111111111111111111111111111111111100"),
		("0000011111111111111111111111111111111111111111111111111111111111"),
		("0011111111111111111111111111111111111111111111111111111111111111"),
		("0011111111111111111111111111111111111111111111111111111111111111"),
		("1111111111111111111111111111111111111111111111111111111111111111"),
		("1111111111111111111111111111111111111111111111111111111111111111"),
		("1111111111111111111111111111111111111111111111111111111111111111"),
		("1111111111111111111111111111111111111111111111111111111111111111"),
		("0011111111111111111111111111111111111111111111111111111111111100"),
		("0011111111111111111111111111111111111111111111111111111111111100"),
		("0000111111111111111111111111111111111111111111111111111111110000"),
		("0000111111111111111111111111111111111111111111111111111111110000"),
		("0000001111111111111111111111111111111111111111111111111111111100"),
		("0000001111111111111111111111111111111111111111111111111111111100"),
		("0000000011111111111111111111111111111111111111111111111111111111"),
		("0000000011111111111111111111111111111111111111111111111111111111"),
		("0000000011111111111111111111111111111111111111111111111111111110"),
		("0000000011111111111111111111111111111111111111111111111111111110"),
		("0000000000111111111111111111111111111111111111111111111111111100"),
		("0000000000111111111111111111111111111111111111111111111111111100"),
		("0000000000000000111111111111111111111111111111111111111111000000"),
		("0000000000000000111111111111111111111111111111111111111111000000"),
		("0000000000000000001111111111111111111111111111111111110000000000"),
		("0000000000000000001111111111111111111111111111111111110000000000"),
		("0000000000000000000000111111111111111111111100000000000000000000"),
		("0000000000000000000000111111111111111111111100000000000000000000")
	);
	
	
	--MATRICE CHE RESTITUISCE IL COLORE DI OGNI PIXEL ASSOCIATO A MARIO
	type nuvola_colori is array (0 to CLOUD_HEIGHT - 1 , 0 to CLOUD_WIDTH - 1) of std_logic_vector(3 downto 0);
	constant cloud_colors : nuvola_colori := (
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"7", x"7", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0"),
		( x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0"),
		( x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0"),
		( x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0"),
		( x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0"),
		( x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0"),
		( x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0"),
		( x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"6", x"6", x"7", x"7", x"6", x"6", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"7", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6", x"6")
	);
	
	
	--MATRICE CHE MI INDICA SE IL PIXEL IDENTIFICA UN ELEMENTO DELLA COLLINA
	type hill_form is array (0 to HILL_HEIGTH - 1 , 0 to HILL_WIDTH - 1) of std_logic;
	constant hill_borders : hill_form := (
		("000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000"),
		("000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000"),
		("000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000"),
		("000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000"),
		("000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000"),
		("000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000"),
		("000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000"),
		("000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000"),
		("000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000"),
		("000000000000000000000000000011111111111111111111111111111111111111110000000000000000000000000000"),
		("000000000000000000000000001111111111111111111111111111111111111111111100000000000000000000000000"),
		("000000000000000000000000001111111111111111111111111111111111111111111100000000000000000000000000"),
		("000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000"),
		("000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000"),
		("000000000000000000000011111111111111111111111111111111111111111111111111110000000000000000000000"),
		("000000000000000000000011111111111111111111111111111111111111111111111111110000000000000000000000"),
		("000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000"),
		("000000000000000000001111111111111111111111111111111111111111111111111111111100000000000000000000"),
		("000000000000000000111111111111111111111111111111111111111111111111111111111111000000000000000000"),
		("000000000000000000111111111111111111111111111111111111111111111111111111111111000000000000000000"),
		("000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000"),
		("000000000000000011111111111111111111111111111111111111111111111111111111111111110000000000000000"),
		("000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000"),
		("000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000"),
		("000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000"),
		("000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000"),
		("000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000"),
		("000000000011111111111111111111111111111111111111111111111111111111111111111111111111110000000000"),
		("000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000"),
		("000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000"),
		("000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000"),
		("000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000"),
		("000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
		("000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
		("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
		("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
		("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111")
	);
	
	
	--
	--MATRICE CHE RESTITUISCE IL COLORE DI OGNI PIXEL ASSOCIATO A MARIO
	type collina_colori is array (0 to HILL_HEIGTH - 1 , 0 to HILL_WIDTH - 1) of std_logic_vector(3 downto 0);
	constant hill_colors : collina_colori := (
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0"),
		( x"0", x"0", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"5", x"0", x"0")
	);
	
	
	--MATRICE CHE MI INDICA SE IL PIXEL IDENTIFICA UN ELEMENTO DEL PAVIMENTO
	type floor_form is array (0 to FLOOR_HEIGTH - 1 , 0 to FLOOR_WIDTH - 1) of std_logic;
	constant floor_borders : floor_form := (
		("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000"),
		("000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000"),
		("000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000"),
		("000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000000110000000000001100000000000011000000000001"),
		("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000"),
		("000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000"),
		("000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000"),
		("000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000"),
		("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("000000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000"),
		("000000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000"),
		("000000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000"),
		("000000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000011000000000")
	);
	
	--MATRICE CHE RESTITUISCE IL COLORE DI OGNI PIXEL ASSOCIATO Al PAVIMENTO
	type floor_colori is array (0 to FLOOR_HEIGTH - 1 , 0 to FLOOR_WIDTH - 1) of std_logic_vector(3 downto 0);
	constant floor_colors : floor_colori := (
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3"),
		( x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3")
	);
	
	--STAR
	--MATRICE CHE MI INDICA SE IL PIXEL IDENTIFICA UN ELEMENTO DELLA STELLA
	type star_form is array (0 to STAR_HEIGHT - 1 , 0 to STAR_WIDTH - 1) of std_logic;
	constant star_borders : star_form := (
		("00000000000011111111000000000000"),
		("00000000000011111111000000000000"),
		("00000000000011111111000000000000"),
		("00000000000011111111000000000000"),
		("00000000000111111111100000000000"),
		("00000000000111111111100000000000"),
		("00000000001111111111110000000000"),
		("00000000001111111111110000000000"),
		("11111111111111111111111111111111"),
		("11111111111111111111111111111111"),
		("11111111111111111111111111111111"),
		("11111111111111111111111111111111"),
		("11111111111111111111111111111111"),
		("11111111111111111111111111111111"),
		("00111111111111111111111111111100"),
		("00111111111111111111111111111100"),
		("00001111111111111111111111110000"),
		("00001111111111111111111111110000"),
		("00000011111111111111111111000000"),
		("00000011111111111111111111000000"),
		("00000011111111111111111111000000"),
		("00000011111111111111111111000000"),
		("00000011111111111111111111000000"),
		("00000011111111111111111111000000"),
		("00000011111111111111111111000000"),
		("00000111111111111111111111100000"),
		("00001111111111111111111111110000"),
		("00001111111111111111111111110000"),
		("00011111111111000011111111111000"),
		("00011111111100000000111111111000"),
		("00111111110000000000011111111100"),
		("00111111110000000000001111111100")
	);
	
	--MATRICE CHE RESTITUISCE IL COLORE DI OGNI PIXEL ASSOCIATO ALLA STELLA
	type star_colori is array (0 to STAR_HEIGHT - 1 , 0 to STAR_WIDTH - 1) of std_logic_vector(3 downto 0);
	constant star_colors : star_colori := (
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0")
	);
	
	type pause_form is array (0 to PAUSE_HEIGHT - 1 , 0 to PAUSE_WIDTH - 1) of std_logic;
	constant pause_borders : pause_form := (
		("11110000000000000000000000000000"),
		("11111100000000000000000000000000"),
		("11001111000000000000000000000000"),
		("11000011110000000000000000000000"),
		("11000000111100000000000000000000"),
		("11000000001111000000000000000000"),
		("11000000000011110000000000000000"),
		("11000000000000111100000000000000"),
		("11000000000000001111000000000000"),
		("11000000000000000011110000000000"),
		("11000000000000000000111100000000"),
		("11000000000000000000001111000000"),
		("11000000000000000000000011110000"),
		("11000000000000000000000000111100"),
		("11000000000000000000000000001111"),
		("11000000000000000000000000000011"),
		("11000000000000000000000000000011"),
		("11000000000000000000000000001111"),
		("11000000000000000000000000111100"),
		("11000000000000000000000011110000"),
		("11000000000000000000001111000000"),
		("11000000000000000000111100000000"),
		("11000000000000000011110000000000"),
		("11000000000000001111000000000000"),
		("11000000000000111100000000000000"),
		("11000000000011110000000000000000"),
		("11000000001111000000000000000000"),
		("11000000111100000000000000000000"),
		("11000011110000000000000000000000"),
		("11001111000000000000000000000000"),
		("11111100000000000000000000000000"),
		("11110000000000000000000000000000")
	);
	
	--MATRICE CHE MI INDICA SE IL PIXEL IDENTIFICA UN ELEMENTO DEI MATTONCINI
	type brick_form is array (0 to 20 - 1 , 0 to 125 - 1) of std_logic;
	constant brick_borders : brick_form := (
		("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("11000000000000110000000000001100000000000011000000000000110000000000000000011000000000000110000000000001100000000000011000011"),
		("11000000000000110000000000001100000000000011000000000000110000000000000000011000000000000110000000000001100000000000011000011"),
		("11000000000000110000000000001100000000000011000000000000110000000000000000011000000000000110000000000001100000000000011000011"),
		("11000000000000110000000000001100000000000011000000000000110000000000000000011000000000000110000000000001100000000000011000011"),
		("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("11000000011000000000011000000000011000000000011000000000011000000000001100000000001100000000001100000000001100000000001100011"),
		("11000000011000000000011000000000011000000000011000000000011000000000001100000000001100000000001100000000001100000000001100011"),
		("11000000011000000000011000000000011000000000011000000000011000000000001100000000001100000000001100000000001100000000001100011"),
		("11000000011000000000011000000000011000000000011000000000011000000000001100000000001100000000001100000000001100000000001100011"),
		("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("11000000000000011000000000011000000000011000000000011000000000000000000000001100000000001100000000001100000000001100000000011"),
		("11000000000000011000000000011000000000011000000000011000000000000000000000001100000000001100000000001100000000001100000000011"),
		("11000000000000011000000000011000000000011000000000011000000000000000000000001100000000001100000000001100000000001100000000011"),
		("11000000000000011000000000011000000000011000000000011000000000000000000000001100000000001100000000001100000000001100000000011"),
		("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
		("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111")
	);
	
	--MATRICE CHE RESTITUISCE IL COLORE DI OGNI PIXEL ASSOCIATO AI MATTONCINI
	type brick_colori is array (0 to BLOCK_HEIGHT - 1 , 0 to BLOCK_WIDTH - 1) of std_logic_vector(3 downto 0);
	constant brick_colors : brick_colori := (
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"3", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0"),
		( x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"0")
	);

	
	type coin_form is array (0 to COIN_HEIGHT - 1 , 0 to COIN_WIDTH - 1) of std_logic;
	constant coin_borders : coin_form := (
		("0000001111000000"),
		("0000011111110000"),
		("0000111111110000"),
		("0001111111111000"),
		("0011111111111100"),
		("0011111111111100"),
		("0011111111111100"),
		("0111111111111110"),
		("0111111111111110"),
		("0111111111111110"),
		("0111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("1111111111111111"),
		("0111111111111111"),
		("0111111111111110"),
		("0111111111111110"),
		("0111111111111110"),
		("0011111111111110"),
		("0011111111111100"),
		("0011111111111100"),
		("0001111111111000"),
		("0000111111110000"),
		("0000011111110000"),
		("0000001111000000")
	);	
	
	type coin_colori is array (0 to COIN_HEIGHT - 1 , 0 to COIN_WIDTH - 1) of std_logic_vector(3 downto 0);
	constant coin_colors : coin_colori := (
		( x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"4", x"4", x"0", x"0", x"0", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"6", x"6", x"6"),
		( x"6", x"6", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"0", x"0", x"4", x"4", x"4", x"4", x"0", x"4", x"4", x"4", x"0", x"0", x"6", x"6"),
		( x"6", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"4", x"4", x"4", x"4", x"0", x"0", x"6"),
		( x"6", x"0", x"0", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"0", x"0", x"6"),
		( x"6", x"0", x"0", x"4", x"4", x"0", x"4", x"4", x"0", x"4", x"0", x"4", x"4", x"0", x"0", x"6"),
		( x"6", x"0", x"0", x"4", x"4", x"0", x"4", x"4", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"0", x"4", x"4", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"0", x"4", x"4", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"0", x"4", x"4", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"0", x"4", x"4", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"4", x"0", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"4", x"0", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"4", x"0", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"4", x"0", x"4", x"4", x"4", x"0", x"0"),
		( x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"4", x"0", x"4", x"4", x"4", x"0", x"0"),
		( x"6", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"4", x"0", x"4", x"4", x"4", x"0", x"0"),
		( x"6", x"0", x"0", x"4", x"4", x"0", x"4", x"4", x"0", x"4", x"0", x"4", x"4", x"0", x"0", x"6"),
		( x"6", x"0", x"0", x"4", x"4", x"4", x"0", x"0", x"0", x"0", x"4", x"4", x"4", x"0", x"0", x"6"),
		( x"6", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"0", x"4", x"4", x"4", x"4", x"0", x"0", x"6"),
		( x"6", x"6", x"0", x"0", x"4", x"4", x"4", x"4", x"0", x"4", x"4", x"4", x"4", x"0", x"0", x"6"),
		( x"6", x"6", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"4", x"4", x"4", x"0", x"0", x"6", x"6"),
		( x"6", x"6", x"6", x"0", x"0", x"0", x"4", x"4", x"4", x"4", x"0", x"0", x"0", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"4", x"4", x"0", x"0", x"0", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6"),
		( x"6", x"6", x"6", x"6", x"6", x"6", x"0", x"0", x"0", x"0", x"6", x"6", x"6", x"6", x"6", x"6")
	);
	
	--SCORE NUMBER
	type number_form is array (0 to CIFRA_HEIGHT - 1 , 0 to CIFRA_WIDTH - 1) of std_logic;
	type double_number_form is array (0 to CIFRA_HEIGHT - 1 , 0 to 2*CIFRA_WIDTH - 1) of std_logic;
	
	constant zero_borders : number_form := (
		("0001111111111000"),
		("0011111111111100"),
		("0110000000000110"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("0110000000000110"),
		("0011111111111100"),
		("0001111111111000")
	);
	
	constant one_borders : number_form := (
		("0000000110000000"),
		("0000001110000000"),
		("0000011110000000"),
		("0000110110000000"),
		("0001100110000000"),
		("0011000110000000"),
		("0110000110000000"),
		("1100000110000000"),
		("1000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0111111111111110"),
		("1111111111111111")
	);	
	
	constant two_borders : number_form := (
		("1111111111111000"),
		("1111111111111100"),
		("0000000000000110"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000110"),
		("0001111111111100"),
		("0011111111111000"),
		("0110000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("0110000000000000"),
		("0011111111111111"),
		("0011111111111111")
		);
	
	constant three_borders : number_form := (
		("1111111111111000"),
		("1111111111111100"),
		("0000000000000110"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000111"),
		("0011111111111110"),
		("0011111111111110"),
		("0000000000000111"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000110"),
		("1111111111111100"),
		("1111111111111000")
	);
	
	constant four_borders : number_form := (
		("0000000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("0110000000000011"),
		("0011111111111111"),
		("0001111111111111"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011")
	);
	
	constant five_borders : number_form := (
		("0001111111111111"),
		("0011111111111111"),
		("0110000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("0110000000000000"),
		("0011111111111000"),
		("0001111111111100"),
		("0000000000000110"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000110"),
		("1111111111111100"),
		("1111111111111000")
	);
	
	constant six_borders : number_form := (
		("0001111111111111"),
		("0011111111111110"),
		("0110000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1100000000000000"),
		("1101111111111000"),
		("1111111111111100"),
		("1110000000000110"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("0110000000000110"),
		("0011111111111100"),
		("0001111111111000")
		);
	
	constant seven_borders : number_form := (
		("1111111111111000"),
		("0111111111111100"),
		("0000000000000110"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011")
		);
	
	constant eight_borders : number_form := (
		("0001111111111000"),
		("0011111111111100"),
		("0110000000000110"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("0110000000000010"),
		("0011111111111100"),
		("0011111111111100"),
		("0110000000000110"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("0100000000000110"),
		("0011111111111100"),
		("0001111111111000")
		);
	
	constant nine_borders : number_form := (
		("0001111111111000"),
		("0011111111111100"),
		("0110000000000110"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("1100000000000011"),
		("0110000000000110"),
		("0011111111111111"),
		("0001111111111111"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000011"),
		("0000000000000110"),
		("1111111111111100"),
		("0111111111111000")
		);
	
	
	constant ten_borders : double_number_form := (
		("00000001100000000001111111111000"),
		("00000011100000000011111111111100"),
		("00000111100000000110000000000110"),
		("00001101100000001100000000000011"),
		("00011001100000001100000000000011"),
		("00110001100000001100000000000011"),
		("01100001100000001100000000000011"),
		("11000001100000001100000000000011"),
		("10000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000001100000000000011"),
		("00000001100000000110000000000110"),
		("00011111111110000011111111111100"),
		("00111111111111000001111111111000")
	);
	
	type t_cifre_array is array(0 to 9) of number_form; -- coordinate type
	constant CIFRE : t_cifre_array := (zero_borders, one_borders, two_borders, three_borders, four_borders, five_borders, six_borders, seven_borders, eight_borders, nine_borders); -- all the blocks are stored here
	
	type x_form is array (0 to X_SCORE_HEIGHT - 1 , 0 to X_SCORE_WIDTH - 1) of std_logic;
	constant x_borders : x_form := (
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0110000000000110"),
		("0110000000000110"),
		("0011000000001100"),
		("0011000000001100"),
		("0001100000011000"),
		("0001100000011000"),
		("0000110000110000"),
		("0000110000110000"),
		("0000011001100000"),
		("0000011001100000"),
		("0000001111000000"),
		("0000001111000000"),
		("0000000110000000"),
		("0000000110000000"),
		("0000001111000000"),
		("0000001111000000"),
		("0000011001100000"),
		("0000011001100000"),
		("0000110000110000"),
		("0000110000110000"),
		("0001100000011000"),
		("0001100000011000"),
		("0011000000001100"),
		("0011000000001100"),
		("0110000000000110"),
		("0110000000000110"),
		("0000000000000000"),
		("0000000000000000")
	);
	
	type eq_form is array (0 to EQUAL_HEIGHT - 1 , 0 to EQUAL_WIDTH - 1) of std_logic;
	constant eq_borders : eq_form := (
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("1111111111111111"),
		("1111111111111111"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("1111111111111111"),
		("1111111111111111"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000"),
		("0000000000000000")
	);
	--FUNCTIONS
	
	--PRENDE IN INGRESSO UN ESADECIMALE E RESTITUISCE LE TRE COMPONENTI RGB
	function get_color(color : in std_logic_vector(3 downto 0))  return matrix_color;
	
end package;

package body vga_package is
	
	function get_color(color : in std_logic_vector(3 downto 0) ) return matrix_color is
	variable RGB : matrix_color;
	begin
			case color is		                  
				when x"0" => RGB(0) := "0000"; RGB(1):="0000"; RGB(2):="0000"; --BLACK
				when x"1" => RGB(0) := "1111"; RGB(1):="1100"; RGB(2):="1101"; --PINK
				when x"2" => RGB(0) := "1111"; RGB(1):="0000"; RGB(2):="0000"; --RED
				when x"3" => RGB(0) := "0111"; RGB(1):="0011"; RGB(2):="0001"; --BROWN LIGHT
				when x"4" => RGB(0) := "1110"; RGB(1):="1101"; RGB(2):="0100"; --YELLOW
				when x"5" => RGB(0) := "0000"; RGB(1):="1111"; RGB(2):="0000"; --GREEN
				when x"6" => RGB(0) := "1111"; RGB(1):="1111"; RGB(2):="1111"; --WHITE
				when x"7" => RGB(0) := "0000"; RGB(1):="1011"; RGB(2):="1111"; --CYAN
				--
				when x"8" => RGB(0) := "0110"; RGB(1):="0001"; RGB(2):="0001"; --BROWN STRONG
				when x"9" => RGB(0) := "0000"; RGB(1):="0000"; RGB(2):="0000"; --BLACK
				when x"A" => RGB(0) := "0000"; RGB(1):="0000"; RGB(2):="0000"; --BLACK
				when x"B" => RGB(0) := "0000"; RGB(1):="0000"; RGB(2):="0000"; --BLACK
				when x"C" => RGB(0) := "0000"; RGB(1):="0000"; RGB(2):="0000"; --BLACK
				when x"D" => RGB(0) := "0000"; RGB(1):="0000"; RGB(2):="0000"; --BLACK
				when x"E" => RGB(0) := "0000"; RGB(1):="0000"; RGB(2):="0000"; --BLACK
				when x"F" => RGB(0) := "0000"; RGB(1):="0000"; RGB(2):="0000"; --BLACK
			end case;

			return RGB;
	 end function;
	
end vga_package;


